module fvtb(input clk, output led);
   blink fvuud (.*);
   always_ff @(posedge clk) begin main: assert(led); wit: cover(led); end
endmodule // fvtb

